//$write work same as $display 
//except it dose not automatically add new line

module write  ;
initial begin
$write("jay shree ram");
$write ("shiyavar ramchandra ki jay ");
$write("satya sanan dharam ki jai ho");
end 
endmodule
