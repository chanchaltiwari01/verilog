module and_gate (c,a,b);
input a,b;
output c;
and (c,a,b);
endmodule
