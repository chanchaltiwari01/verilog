//$display use to display of value and statement
//it is execute at active region 
//execute in 0 simulaton time/ insert new line by default 
module display ;
initial begin
$display("jay shree ram");
$display ("shiyavar ramchandra ki jay ");
$display("satya sanan dharam ki jai ho");
end 
endmodule
